module raymath

#flag -I @VMODROOT/raymath/
#flag @VMODROOT/raymath/raymath.h
#include "raymath.h"
