module raygui

#flag -I @VMODROOT/raygui/
#flag @VMODROOT/raygui/raygui.h
#define RAYGUI_IMPLEMENTATION
#include "raygui.h"
