module raymath

#flag -I @VMODROOT/raymath/
#include "raymath.h"
