module raygui

#flag -I @VMODROOT/raygui/
#define RAYGUI_IMPLEMENTATION
#include "raygui.h"
